module multiplier_toplevel
(

    input   logic           Clk,        // 50MHz clock is only used to get timing estimate data
    input   logic           Reset,      // From push-button 0.  Remember the button is active low (0 when pressed)
    input   logic           Run,        // From push-button 3.
    input   logic           ClearA_LoadB,         // From slider switches
	 input 	logic	[7:0]		 S,
	 
	 output  logic [6:0]  	 AhexL,				// Hex drivers display both inputs to the adder.
									 AhexU,
									 BhexL,
									 BhexU,
	 output  logic [7:0] 	 Aval, 
									 Bval,
	 output  logic 			 X);

// Need module that describes control 
    logic          Clr_A;      // From push-button 1
	 logic          Shift;      // From push-button 1
	 logic          Add;      // From push-button 1
	 logic          Sub;      // From push-button 1
	 logic[7:0]     A;  // Shift register A
	 logic[7:0]     B;  // Shift register B
	 logic[8:0]     Aout;  // Shift register A
	 logic 			 Xout;  // Sign extension bit 
	 logic 			 LSB;
	 
	 assign LSB = B[0];
	 
	 
	ninebit_adder 		addition_unit (
							.A(A),
							.S(S^Sub),
							.M(Sub),
							.AxS(Aout),
							.X(Xout));
	reg_8					register_unitA  ( 		// come back to these imputs
							.Clk(Clk), 
							.Reset(Reset), 
							.Shift_In(A[7]), 
							.Load(ClearA_LoadB), 
							.Shift_En(Shift),
							.D(S));
	reg_8					register_unitB  (
							.Clk(Clk), 
							.Reset(Reset), 
							.Shift_In(B[7]), 
							.Load(ClearA_LoadB), 
							.Shift_En(Shift),
							.D(S));
	control_logic		control_unit (
							.Add(Add),
							.Sub(Sub),
							.Shift(Shift),
							.Clr_A(Clr_A)
							);
	 
	 always_ff @(posedge Clk) begin
        
        if (Clr_A) begin
            // if clear var is high, clear A
            A <= 8'h000;
            X <= 1'b0;
        end else if (!Reset) begin
            // if reset is pressed, clear the adder's input registers
            A <= 8'h000;
            B <= 8'h000;
            X <= 1'b0;
        end else if (!ClearA_LoadB) begin
            // if reset is pressed, clear the adder's input registers
            A <= 8'h000;
            B <= S;
            X <= 1'b0;
        end else if (Add && LSB) begin
				A <= Aout[7:0]; 
				X <= Xout;
		  end else if (Shift) begin
				B = B	>> 1;
				B[7] = A[0];
				A = A >>> 1;
				A[7] = X;
		  end 
	 end

//	  sync button_sync[3:0] (Clk, {~Reset, ~Run, ClearA_LoadB}, {Reset_SH, Run_SH, LoadB_SH, Execute_SH});
//	  sync Din_sync[7:0] (Clk, Din, Din_S);
//	  sync F_sync[2:0] (Clk, F, F_S);
//	  sync R_sync[1:0] (Clk, R, R_S);
	

endmodule