module datapath ();


//Todo:
/* -instantiate PC, Address ALU, BUS, MAR, MDR, IR, Reg_file, ALU, CC, testbench lol */



endmodule 

