module PC (); //Program Counter Register, stores address of next instruction


endmodule 

module Address_ALU (input offset, //ALU near PC that computes the next PC value based on current instruction
						  input offset_flag,
						  output address); //flag whether should comput using offet or just be PC + 1
						  
						  
endmodule 

module BUS ();


endmodule

module MAR ();


endmodule

module MDR ();


endmodule

module IR ();


endmodule 

module Reg_file ();


endmodule 

module ALU ();


endmodule 

module CC ();


endmodule 